`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// AY1718 Sem 1 EE2020 Project
// Project Name: Audio Effects
// Module Name: AUDIO_FX_TOP
// Team No.: 
// Student Names: 
// Matric No.:
// Description: 
// 
// Work Distribution:
//////////////////////////////////////////////////////////////////////////////////

module AUDIO_FX_TOP(
    input CLK,            // 100MHz FPGA clock
    input [1:0] caseSwitch, //switch between the 4 cases
    input [10:0] sw, //switch for music instrument
    input [1:0] swD, //switch for delay
    
    input reset,    //buttons
    input left, right,
    
    
    input  J_MIC3_Pin3,   // PmodMIC3 audio input data (serial)
    output J_MIC3_Pin1,   // PmodMIC3 chip select, 20kHz sampling clock
    output J_MIC3_Pin4,   // PmodMIC3 serial clock (generated by module SPI.v)
     
    output J_DA2_Pin1,    // PmodDA2 sampling clock (generated by module DA2RefComp.vhd)
    output J_DA2_Pin2,    // PmodDA2 Data_A, 12-bit speaker output (generated by module DA2RefComp.vhd)
    output J_DA2_Pin3,    // PmodDA2 Data_B, not used (generated by module DA2RefComp.vhd)
    output J_DA2_Pin4,    // PmodDA2 serial clock, 50MHz clock
    
    output reg Hsync, Vsync,
    output [11:0] rgb,
    
    // Seven segment display outputs
    output  [3:0] an,
    output  [6:0] seg,
    output  dp,
    // Seven segment display outputs
    output reg [11:0] led
    );

    //////////////////////////////////////////////////////////////////////////////////
    // Clock Divider Module: Generate necessary clocks from 100MHz FPGA CLK
    // Please create the clock divider module and instantiate it here.
      wire clk_20k;
      wire clk_50M;
      
      get_clock_20k f1(CLK, clk_20k);
      get_clock_50M f2(CLK, clk_50M);
  
     //////////////////////////////////////////////////////////////////////////////////
     //SPI Module: Converting serial data into a 12-bit parallel register
     //Do not change the codes in this area
     //led to observe the effects of MIC_in
       wire [11:0]MIC_in;
       SPI u1 (CLK, clk_20k, J_MIC3_Pin3, J_MIC3_Pin1, J_MIC3_Pin4, MIC_in);
       
       always @ (posedge clk_20k) begin
           led = MIC_in;
       end


    /////////////////////////////////////////////////////////////////////////////////////
    // Real-time Audio Effect Features
    // Please create modules to implement different features and instantiate them here   
     reg [11:0] speaker_out;
     wire [11:0] music;
     wire [11:0] extra_feature;
     wire [11:0] delay;
     
    // wire [6:0] display1, display2;
     wire [3:0] score;
     wire Hsync_temp, Vsync_temp;
     
     A_delay a1(MIC_in, swD, clk_20k, delay);
    
     music_instrument ms(CLK, sw[10:7], sw[6:0], music);  
     vga_pong vp(CLK, reset, left, right, Hsync_temp, Vsync_temp, rgb, extra_feature);
     
     //////////EXTRA FEATURE///////////////////////////
     //////////1. Seven Segment Display//////////////////
     //////////2. VGA PONG GAME + 7 SEGMENT DISPLAY
 
     SSD seg_display (CLK, caseSwitch, sw, swD, an, seg, dp);

     /////////////////////////////////////////////////////////////////////////////
     // assign speaker_out to any of the 4 cases by controlling to switch
    /////////////////////////////////////////////////////////////////////////////////////
    //DAC Module: Digital-to-Analog Conversion
    //Do not change the codes in this area       
    always @ (caseSwitch) begin
        case (caseSwitch)
            2'b00 : speaker_out <= MIC_in;
            2'b01 : speaker_out <= delay;
            2'b10 : speaker_out <= music;
            2'b11 : begin speaker_out <= extra_feature; Hsync <= Hsync_temp; Vsync <= Vsync_temp; end
        endcase
    end
             

     DA2RefComp u2(clk_50M, clk_20k, speaker_out, ,1'b0, J_DA2_Pin2, J_DA2_Pin3, J_DA2_Pin4, J_DA2_Pin1,);
        
  //////////////////////////////////////////////////////////////////////////////////

endmodule
